module single_cycle_mips (
    input logic clk, // clock signal
    input logic rst_n // active-low reset signal used for initialization
);
    
endmodule